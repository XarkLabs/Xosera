// xosera_tb.sv
//
// vim: set et ts=4 sw=4
//
// Copyright (c) 2020 Xark - https://hackaday.io/Xark
//
// See top-level LICENSE file for license information. (Hint: MIT)
//
//`default_nettype none    // mandatory for Verilog sanity
//`timescale 1ns/1ps

`include "xosera_pkg.sv"

`default_nettype none               // mandatory for Verilog sanity
`timescale 1ns/1ps                  // mandatory to shut up Icarus Verilog

module xosera_def_files();

import xv::*;

/* verilator lint_off UNUSED */

typedef enum {
    lang_c,
    lang_asm
} lang_t;

lang_t lang;
integer file;

initial begin
            $display("Xosera - dumping definitions");

            write_defs_lang(lang_c);
            write_defs_lang(lang_asm);

end

task write_defs_lang(
        lang_t  l
    );
    begin
        lang = l;
        file = -1;
        case (lang)
            lang_c:     begin
                file = $fopen("sim/logs/xosera_test_defs.h", "w");
                write_comment("xosera_defs.h");
            end
            lang_asm:   begin
                    file = $fopen("sim/logs/xosera_test_defs.inc", "w");
                    write_comment("xosera_defs.inc");
            end
            default:
                $error("bad lang");
        endcase
            write_comment("NOTE: Do not edit, this is auto-generated by `make def_files` using");
            write_comment("      xosera_pkg.sv file as the one source of truth.");
            write_blank();
            write_comment("Xosera main registers (16-bit, directly accessible)");
            write_reg_def(0, "system control register with a really really long comment");
            write_reg_def(1, "system interrupt control register with a really really long comment");
        $fclose(file);
        file = -1;
    end
endtask

task write_blank(
    );
    begin
        $fwrite(file, "\n");
    end
endtask

task write_comment(
        input logic [128*8-1:0]  comment
    );
    begin
        case (lang)
            lang_c:
                $fwrite(file, "// %-s\n", comment);
            lang_asm:
                $fwrite(file, "; %-s\n", comment);
            default:
                $error("bad lang");
        endcase
    end
endtask

task write_reg_def(
        input logic [7:0]   num,
        input logic [128*8-1:0]  comment
    );
    begin
        case (lang)
            lang_c:
                $fwrite(file, "#define     %-16s    0x%02x    // %-s\n", regname(4'(num)), num, comment);
            lang_asm:
                $fwrite(file, "%-16s    =   $%02x     ; %-s\n", regname(4'(num)), num, comment);
            default:
                $error("bad lang");
        endcase
    end
endtask

function automatic logic [63:0] regname(
        input logic [3:0] num
    );
    begin
        case (num)
            4'h0: regname = "XR_ADDR ";
            4'h1: regname = "XR_DATA ";
            4'h2: regname = "RD_INCR ";
            4'h3: regname = "RD_ADDR ";
            4'h4: regname = "WR_INCR ";
            4'h5: regname = "WR_ADDR ";
            4'h6: regname = "DATA    ";
            4'h7: regname = "DATA2   ";
            4'h8: regname = "SYS_CTRL";
            4'h9: regname = "TIMER   ";
            4'hA: regname = "UNUSED_A";
            4'hB: regname = "UNUSED_B";
            4'hC: regname = "RW_INCR ";
            4'hD: regname = "RW_ADDR ";
            4'hE: regname = "RW_DATA ";
            4'hF: regname = "RW_DATA2";
            default: regname = "????????";
        endcase
    end
endfunction

endmodule

`default_nettype wire               // restore default
